// *****************************************************
// AVR address constants (localparams)
//  for registers used by Xcelerator Blocks (XBs) 
// *****************************************************

localparam PAD0_ADDR  = 8'hE0;
localparam PAD1_ADDR  = 8'hE1;
localparam PNGCR_ADDR = 8'hE2;

